module int32u(
    input int32_opc,
    input int32_a,
    input int32_b,
    output int32_y,
    input int32_iv,
    input int32_or,
    output int32_ov,
    output int32_ir
)
endmodule