module uint32Unit(
    input uint32_opc,
    input uint32_a,
    input uint32_b,
    output uint32_y,
    input uint32_iv,
    input uint32_or,
    output uint32_ov,
    output uint32_ir
)
endmodule